`include "defines.v"
`include "start_detect_tb.v"
`include "start_detec_tester.v"


module start_detect_tb;
   


endmodule // start_detect_tb

