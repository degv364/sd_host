`include "defines.v"

module delayer(input clk,
	       input [31:0] data_in,
	       output [31:0] data_out);
   
   reg [31:0] 		     memory;
   
   always @(posedge clk) begin


      endmodule // delayer

   
