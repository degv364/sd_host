`include "defines.v"


module start_detect_tester();



endmodule // start_detect_tester
